LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY setting IS
    PORT (
        sel : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        output : OUT STD_LOGIC_VECTOR(50 DOWNTO 0)
    );
END setting;

ARCHITECTURE RTL OF setting IS
BEGIN
    PROCESS (sel)
    BEGIN
        CASE sel IS
            WHEN "0000" =>
                output <= "000000000000000000000000000100000000000000000000001";
            WHEN "0001" =>
                output <= "000000000000000000000000010000000000000000000000001";
            WHEN "0010" =>
                output <= "000000000000000000000000100000000000000000000000001";
            WHEN "0011" =>
                output <= "000000000000000000000100000000000000000000000000001";
            WHEN "0100" =>
                output <= "000000000000000001000000000000000000000000000000001";
            WHEN "0101" =>
                output <= "000000000000000100000000000000000000000000000000001";
            WHEN "0110" =>
                output <= "000000000001000000000000000000000000000000000000001";
            WHEN "0111" =>
                output <= "001000000000000000000000000000001000000000000000001";
            WHEN "1000" =>
                output <= "000000000000000000000000000000100000000000000000001";
            WHEN "1001" =>
                output <= "000000000000000010000000000000000000000000000000001";
            WHEN "1010" =>
                output <= "000000000000000000000000000000000000000000010000001";
            WHEN "1011" =>
                output <= "000000000000000000000000000000000100000000000000001";
            WHEN "1100" =>
                output <= "000000000000000000000000000000000000000000000010001";
            WHEN "1101" =>
                output <= "000000000000000000000000000000000000000000000100001";
            WHEN "1110" =>
                output <= "000000000000000000000000000000000000000000000000011";
            WHEN "1111" =>
                output <= "000000000000000000000000000000000000000000000000010";

                -- Default case: if none of the above selectors match
            WHEN OTHERS =>
                output <= "000000000000000000000000000000000000000000000000000";
        END CASE;
    END PROCESS;
END RTL;